FWD,29052016:09:01,10.56| FWD,29052016:10:53,11.23| FWD,29052016:15:40,23.20
SPOT,29052016:09:04,11.56| FWD,29052016:11:45,11.23| SPOT,29052016:12:30,23.20
FWD,29052016:08:01,10.56| SPOT,29052016:12:30,11.23| FWD,29052016:13:20,23.20| FWD,29052016:14:340,56.00
FWD,29052016:08:01,10.56| SPOT,29052016:12:30,11.23| FWD,29052016:13:20,23.20
